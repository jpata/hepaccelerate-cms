jobfiles/dy_2017_142.json
jobfiles/ttjets_sl_2018_29.json
jobfiles/data_2018_452.json
jobfiles/data_2017_74.json
jobfiles/data_2017_41.json
