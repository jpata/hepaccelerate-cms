jobfiles/wz_2l2q_2016_0.json
jobfiles/data_2016_344.json
jobfiles/data_2016_286.json
jobfiles/data_2018_84.json
jobfiles/st_tw_top_2017_7.json
